`timescale 1ns / 1ps
`default_nettype none

module crossp_tb();
    logic clk_in;

    logic [31:0] vector1_x;
    logic [31:0] vector1_y;
    logic [31:0] vector1_z;

    logic [31:0] vector2_x;
    logic [31:0] vector2_y;
    logic [31:0] vector2_z;

    logic [31:0] cross_vec_x;
    logic [31:0] cross_vec_y;
    logic [31:0] cross_vec_z;

    logic data_valid_in;
    logic data_valid_out;
    logic vectors_ready;

    cp_wrapper uut(
      .clk_in(clk_in),
      .valid_in(data_valid_in),
      .vec_ax(vector1_x), 
      .vec_ay(vector1_y), 
      .vec_az(vector1_z), 
      .vec_bx(vector2_x),
      .vec_by(vector2_y),
      .vec_bz(vector2_z),
      .vec_ready(vectors_ready),
      .value_out_x(cross_vec_x),
      .value_out_y(cross_vec_y),
      .value_out_z(cross_vec_z),
      .valid_out(data_valid_out),
      .cross_product_ready(1'b1)
    );

    always begin
      #5;  //every 5 ns switch...so period of clock is 10 ns...100 MHz clock
      clk_in = !clk_in;
    end

    //https://www.h-schmidt.net/FloatConverter/IEEE754.html
    
    initial begin
      $dumpfile("crossp_tb.vcd"); //file to store value change dump (vcd)
      $dumpvars(0,crossp_tb);
      $display("Starting Sim"); //print nice message at start
      clk_in = 0;
      #10;
      vector1_x = 32'h4080_0000; // 4 in floating point notation
      vector1_y = 32'h4110_0000; // 9 in floating point notation
      vector1_z = 32'h0;
      vector2_x = 32'h3f80_0000; // 1 in floating point notation
      vector2_y = 32'h0;
      vector2_z = 32'h0;
      data_valid_in = 1;
      #10;
      data_valid_in = 0;
      #2000;
      $finish;
    end
endmodule

`default_nettype wire